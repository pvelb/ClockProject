module TestMudule1

input wire port_a,
output wire port_b,

port_b=port_a;

endmodule